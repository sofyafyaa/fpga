module dec_3x8(input en,
					input [3:0] in, 	 
					output reg [15:0] out);
				
	always @(en or in) begin
		out = en ? 1 << in: 0;
	end
endmodule